module main

import hello_world

fn main() {
	println(hello_world.hello_world())
}
