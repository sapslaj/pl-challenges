module hello_world

pub fn hello_world() string {
	return 'hello world'
}
